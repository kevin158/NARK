module _NOT(input logic X, output logic Y);
	assign Y = ~X;
endmodule 