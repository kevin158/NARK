module SIXTY_FOUR_N_BITS_INPUTS_SIX_BITS_SELECT_MUX_MODULE #(parameter BITS = 32) (DATA, SELECT, OUT);

	input logic [63:0][BITS-1:0] DATA;
	input logic [5:0] SELECT;
	output logic [BITS-1:0] OUT;
	logic [BITS-1:0] W_FIRST_MUX, W_SECOND_MUX;
	
	THIRTY_TWO_N_BITS_INPUTS_FIVE_BITS_SELECT_MUX_MODULE #(BITS)
		FIRST_MUX (DATA[31:0], SELECT[4:0], W_FIRST_MUX),
		SECOND_MUX (DATA[63:32], SELECT[4:0], W_SECOND_MUX);
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS)
		THIRD_MUX (W_FIRST_MUX, W_SECOND_MUX, SELECT[5], OUT);
	
endmodule 