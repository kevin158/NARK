module SIX_BITS_SELECT_SIXTY_FOUR_DEMUX_MODULE (IN, SELECT, OUT);
	
	input  logic 		  IN;
	input  logic [5:0]  SELECT;
	output logic [63:0] OUT;
	logic        [15:0]  W_IN;
	
	FOUR_BITS_SELECT_SIXTEEN_DEMUX_MODULE 
		MAIN_DEMUX (IN, SELECT[5:2], W_IN);
	FOUR_BITS_SELECT_SIXTEEN_DEMUX_MODULE
		DEMUX_1  (W_IN[0],  SELECT[1:0], OUT[3:0]),
		DEMUX_2  (W_IN[1],  SELECT[1:0], OUT[7:4]),
		DEMUX_3  (W_IN[2],  SELECT[1:0], OUT[11:8]),
		DEMUX_4  (W_IN[3],  SELECT[1:0], OUT[15:12]),
		DEMUX_5  (W_IN[4],  SELECT[1:0], OUT[19:16]),
		DEMUX_6  (W_IN[5],  SELECT[1:0], OUT[23:20]),
		DEMUX_7  (W_IN[6],  SELECT[1:0], OUT[27:24]),
		DEMUX_8  (W_IN[7],  SELECT[1:0], OUT[31:28]),
		DEMUX_9  (W_IN[8],  SELECT[1:0], OUT[35:32]),
		DEMUX_10 (W_IN[9],  SELECT[1:0], OUT[39:36]),
		DEMUX_11 (W_IN[10], SELECT[1:0], OUT[43:40]),
		DEMUX_12 (W_IN[11], SELECT[1:0], OUT[47:44]),
		DEMUX_13 (W_IN[12], SELECT[1:0], OUT[51:48]),
		DEMUX_14 (W_IN[13], SELECT[1:0], OUT[55:52]),
		DEMUX_15 (W_IN[14], SELECT[1:0], OUT[59:56]),
		DEMUX_16 (W_IN[15], SELECT[1:0], OUT[63:60]);
		
endmodule 