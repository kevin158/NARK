module _OR(input logic X,Y, output logic Z);
	assign Z = X | Y;
endmodule