module FIVE_BITS_SELECT_THIRTY_TWO_DEMUX_MODULE (IN, SELECT, OUT);
	
	input  logic 		  IN;
	input  logic [4:0]  SELECT;
	output logic [31:0] OUT;
	logic        [15:0]  W_IN;
	
	FOUR_BITS_SELECT_SIXTEEN_DEMUX_MODULE 
		MAIN_DEMUX (IN, SELECT[4:1], W_IN);
	ONE_BITS_SELECT_TWO_DEMUX_MODULE
		DEMUX_1  (W_IN[0],  SELECT[0], OUT[1:0]),
		DEMUX_2  (W_IN[1],  SELECT[0], OUT[3:2]),
		DEMUX_3  (W_IN[2],  SELECT[0], OUT[5:4]),
		DEMUX_4  (W_IN[3],  SELECT[0], OUT[7:6]),
		DEMUX_5  (W_IN[4],  SELECT[0], OUT[9:8]),
		DEMUX_6  (W_IN[5],  SELECT[0], OUT[11:10]),
		DEMUX_7  (W_IN[6],  SELECT[0], OUT[13:12]),
		DEMUX_8  (W_IN[7],  SELECT[0], OUT[15:14]),
		DEMUX_9  (W_IN[8],  SELECT[0], OUT[17:16]),
		DEMUX_10 (W_IN[9],  SELECT[0], OUT[19:18]),
		DEMUX_11 (W_IN[10], SELECT[0], OUT[21:20]),
		DEMUX_12 (W_IN[11], SELECT[0], OUT[23:22]),
		DEMUX_13 (W_IN[12], SELECT[0], OUT[25:24]),
		DEMUX_14 (W_IN[13], SELECT[0], OUT[27:26]),
		DEMUX_15 (W_IN[14], SELECT[0], OUT[29:28]),
		DEMUX_16 (W_IN[15], SELECT[0], OUT[31:30]);
		
endmodule 