module REGISTER_FILE_MODULE #(parameter BITS = 24) (CLK, RST, ADDRS_RN, ADDRS_RM, ADDRS_RD, WRT_DATA, R15_DATA, WRT_ENA, RN_DATA, RM_DATA);
	
	input logic             CLK, RST, WRT_ENA;
	input logic  [3:0]      ADDRS_RN, ADDRS_RM, ADDRS_RD;
	input logic  [BITS-1:0] WRT_DATA, R15_DATA;
	output logic [BITS-1:0] RN_DATA, RM_DATA;
	
	logic [15:0] 		      DEMUX_WRITE;
	logic [15:0] [BITS-1:0] REGISTER_DATA;
	logic [BITS-1:0]        WRT_DATA_R15_MUX;
	
	logic                   W_WRITE_R12, W_WRITE_R14, Cout, W_AND_ENA_MUX;
	logic [BITS-1:0]        W_SHIFT_R12, 
	                        W_ADD_R14, 
							      W_WRITE_DATA_R12, 
									W_WRITE_DATA_R14, 
									REGISTER_DATA_R12, 
									REGISTER_DATA_R13, 
									REGISTER_DATA_R14,
									SHIFTED_R12,
									MULTIPLIED_R13,
									ADDED_R14,
									W_ASR_R12,
									W_ASR_R13,
									W_ADD_R13_MUX;
	
	FOUR_BITS_SELECT_SIXTEEN_DEMUX_MODULE 
		FBSSDM (WRT_ENA, ADDRS_RD, DEMUX_WRITE);
	
	REGISTER_MODULE #(BITS,1'b0)
		R0  (CLK, RST, DEMUX_WRITE[0],  WRT_DATA,  		  REGISTER_DATA[0]),
		R1  (CLK, RST, DEMUX_WRITE[1],  WRT_DATA, 		  REGISTER_DATA[1]),
		R2  (CLK, RST, DEMUX_WRITE[2],  WRT_DATA, 		  REGISTER_DATA[2]),
		R3  (CLK, RST, DEMUX_WRITE[3],  WRT_DATA, 		  REGISTER_DATA[3]),
		R4  (CLK, RST, DEMUX_WRITE[4],  WRT_DATA, 		  REGISTER_DATA[4]),
		R5  (CLK, RST, DEMUX_WRITE[5],  WRT_DATA,         REGISTER_DATA[5]),
		R6  (CLK, RST, DEMUX_WRITE[6],  WRT_DATA,         REGISTER_DATA[6]),
		R7  (CLK, RST, DEMUX_WRITE[7],  WRT_DATA,         REGISTER_DATA[7]),
		R8  (CLK, RST, DEMUX_WRITE[8],  WRT_DATA,         REGISTER_DATA[8]),
		R9  (CLK, RST, DEMUX_WRITE[9],  WRT_DATA,         REGISTER_DATA[9]),
		R10 (CLK, RST, DEMUX_WRITE[10], WRT_DATA,         REGISTER_DATA[10]),
		R11 (CLK, RST, DEMUX_WRITE[11], WRT_DATA,         REGISTER_DATA[11]),
		R12 (~CLK, RST, W_WRITE_R12,     W_WRITE_DATA_R12, REGISTER_DATA[12]),
		R13 (CLK, RST, DEMUX_WRITE[13], WRT_DATA,         REGISTER_DATA[13]),
		R14 (~CLK,RST, W_WRITE_R14,     W_WRITE_DATA_R14, REGISTER_DATA[14]),
		R15 (CLK, RST, 1'b1,            WRT_DATA_R15_MUX, REGISTER_DATA[15]); 
	 
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS) 
		NBOSMM (R15_DATA, WRT_DATA, DEMUX_WRITE[15], WRT_DATA_R15_MUX); 
				
	SIXTEEN_N_BITS_INPUTS_FOUR_BITS_SELECT_MUX_MODULE #(BITS) 
		RN_SNBIFBSMM (REGISTER_DATA, ADDRS_RN, RN_DATA),
		RM_SNBIFBSMM (REGISTER_DATA, ADDRS_RM, RM_DATA);

//--------------------------------------------------------------------------------------------------------------	
//Specific purpose register hardware for kernel improvement (R12 =  Kernel row, R14 = Processed pixel)
//--------------------------------------------------------------------------------------------------------------
	
	ONE_BIT_MUX_MODULE
		WRT_R12_MUX (DEMUX_WRITE[13], DEMUX_WRITE[12], DEMUX_WRITE[12], W_WRITE_R12),
		WRT_R14_MUX (DEMUX_WRITE[13], DEMUX_WRITE[14], DEMUX_WRITE[14], W_WRITE_R14);
	
	assign REGISTER_DATA_R12 = REGISTER_DATA[12];
	assign REGISTER_DATA_R13 = REGISTER_DATA[13];
	assign REGISTER_DATA_R14 = REGISTER_DATA[14];
	
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS)
		DATA_R12_MUX (SHIFTED_R12,    WRT_DATA,  DEMUX_WRITE[12], W_WRITE_DATA_R12),
		DATA_R14_MUX (ADDED_R14,      WRT_DATA,  DEMUX_WRITE[14], W_WRITE_DATA_R14),
		DATA_R13_MUX (MULTIPLIED_R13, W_ASR_R13, ~ W_AND_ENA_MUX,   W_ADD_R13_MUX);
	
	N_BITS_LOGIC_SHIFT_LEFT #(BITS)
		LSR_R12 (REGISTER_DATA_R12, BITS/3, SHIFTED_R12);
	 
	N_BITS_ARITMETIC_SHIFT_RIGHT #(BITS)
		ASR_R12 (REGISTER_DATA_R12, BITS-(BITS/3), W_ASR_R12),
		ASR_R13 (REGISTER_DATA_R13, 24'd3,         W_ASR_R13);
	
	N_BITS_MULTIPLIER #(BITS)
		MUL_R13 (REGISTER_DATA_R13, W_ASR_R12, MULTIPLIED_R13);
	 
	ADDER_MODULE #(BITS)
		ADD_R14 (W_ADD_R13_MUX, REGISTER_DATA_R14, 1'b0, ADDED_R14, Cout);
	
	N_INPUTS_OR #(BITS) 
		SHIFT_NIA (REGISTER_DATA_R12, W_AND_ENA_MUX);
 
endmodule 