module _AND(input logic X,Y, output logic Z);
	assign Z = X & Y;
endmodule