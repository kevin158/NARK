module FOUR_N_BITS_INPUTS_TWO_BITS_SELECT_MUX_MODULE #(parameter BITS = 32) (DATA, SELECT, OUT);

	input logic [3:0][BITS-1:0] DATA;
	input logic [1:0] SELECT;
	output logic [BITS-1:0] OUT;
	logic [BITS-1:0] W_FIRST_MUX, W_SECOND_MUX;
	
	N_BITS_ONE_SELECT_MUX_MODULE #(BITS)
		FIRST_MUX (DATA[0], DATA[1], SELECT[0], W_FIRST_MUX),
		SECOND_MUX (DATA[2], DATA[3], SELECT[0], W_SECOND_MUX),
		THIRD_MUX (W_FIRST_MUX, W_SECOND_MUX, SELECT[1], OUT);
	
endmodule 